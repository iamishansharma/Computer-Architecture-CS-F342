module instructionmemory(Inst, PC, clk);

	input[31:0] PC;
	input clk;
	output[31:0] Inst;
	reg [31:0] memory [0:31];
	reg [31:0] Inst;
    integer addr;

    initial 
    begin
	    memory[0] = 32'b00000000000000000000000000000000;  // nop
	    memory[1] = 32'b00000000000000000000000000000000;  // nop
	    memory[2] = 32'b00000000000000000000000000000000;  // nop
	    memory[3] = 32'b00000000000000000000000000000000;  // nop
	    memory[4] = 32'b00000000000000000000000000000000;  // nop
	    memory[5] = 32'b00000000000000000000000000000000;  // nop
	    memory[6] = 32'b00000000000000000000000000000000;  // nop
	    memory[7] = 32'b00000000000000000000000000000000;  // nop
	    memory[8] = 32'b00000000000000000000000000000000;  // nop
	    memory[9] = 32'b00000000000000000000000000000000;  // nop
	    memory[10]= 32'b00000000000000000000000000000000;  // nop
	    memory[11]= 32'b00000000000000000000000000000000;  // nop
	    memory[12]= 32'b00000000000000000000000000000000;  // nop
	    memory[13]= 32'b00000000000000000000000000000000;  // nop
	    memory[14]= 32'b00000000000000000000000000000000;  // nop
	    memory[15]= 32'b00000000000000000000000000000000;  // nop
	    memory[16]= 32'b00000000000000000000000000000000;  // nop
	    memory[17]= 32'b00000000000000000000000000000000;  // nop
	    memory[18]= 32'b00000000000000000000000000000000;  // nop 
	    memory[19]= 32'b00000000000000000000000000000000;  // nop
	    memory[20]= 32'b00000000000000000000000000000000;  // nop
	    memory[21]= 32'b00000000000000000000000000000000;  // nop
	    memory[22]= 32'b00000000000000000000000000000000;  // nop
	    memory[23]= 32'b00000000000000000000000000000000;  // nop
	    memory[24]= 32'b00000000000000000000000000000000;  // nop
	    memory[25]= 32'b00000000000000000000000000000000;  // nop
	    memory[26]= 32'b00000000000000000000000000000000;  // nop
	    memory[27]= 32'b00000000000000000000000000000000;  // nop
	    memory[28]= 32'b00000000000000000000000000000000;  // nop 
	    memory[29]= 32'b00000000000000000000000000000000;  // nop
	    memory[30]= 32'b00000000000000000000000000000000;  // nop
	    memory[31]= 32'b00000000000000000000000000000000;  // nop
  	end

  	always @(posedge clk) 
  	begin
	    addr = PC[31:0];
	    Inst = memory[addr/4];
	end

endmodule